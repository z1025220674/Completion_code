

//function：generate row vector of matrix
module csc_stor #(
    MAT_RANK    =   256
) (
    input                                       clk,
    input                                       rst_n,

    input               
    input               [31     : 0]            s_val_i,
    input               [31     : 0]            s_val_r,
    input               [31     : 0]            a0_val_i,
    input               [31     : 0]            a0_val_r,
    input               [31     : 0]            a1_val_i,
    input               [31     : 0]            a1_val_r,
    input                                       val_vld

);
    



    
endmodule