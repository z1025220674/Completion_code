module sparse_mat #(
    
) (
    
);
    
endmodule