//===================================
//date:2023/1/9
//function:generate sparse matrix and store by csc format
//email:1025220674@qq.com
//vivado2018.3
//===================================
module mat_csc #(
    parameter  = ,
) (
    
);
    
endmodule